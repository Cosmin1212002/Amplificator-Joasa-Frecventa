** Profile: "SCHEMATIC1-Simulari"  [ C:\Users\Fierea Cosmin\Desktop\P1_2024_431D_Fierea_Cosmin-Andrei_AAF_N15_OrCAD\Schematics\p1-pspicefiles\schematic1\simulari.sim ] 

** Creating circuit file "Simulari.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Users\Fierea Cosmin\AppData\Roaming\SPB_16.6\cdssetup\OrCAD_PSpice\17.2.0\PSpice.ini file:
.lib "nomd.lib" 

*Analysis directives: 
.TRAN  0 3m 0 1u 
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
